module inverter(
    input a,
    output a_invert
);

    assign a_invert = invert;

endmodule